`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    06:38:31 04/14/2015 
// Design Name: 
// Module Name:    map 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module map_generator(clk_vga, reset, CurrentX, CurrentY, HBlank, VBlank, playerColor, mapData,
							mapX, mapY
    );

	input [9:0]CurrentX;
	input [8:0]CurrentY;
	input [7:0]playerColor;
	input [3:0]mapX;
	input [3:0]mapY;
	input clk_vga;
	input reset;
	input HBlank;
	input VBlank;
	
	output [7:0]mapData;
	
	reg [7:0]mColor;
	
	//Rooms
	wire [7:0]startCastle;
	wire [7:0]hallwayTop;
	wire [7:0] hallwayRight;
	wire [7:0] blackKeyRoom;
	wire [7:0] hallwayLeft;
	
	//Each map layout is split into its own module for readability
	StartCastle StartCastle(
		.clk_vga(clk_vga),
		.CurrentX(CurrentX),
		.CurrentY(CurrentY),
		.mapData(startCastle),
		.wall(playerColor)
	);
	
	HallwayTop HallwayTop(
		.clk_vga(clk_vga),
		.CurrentX(CurrentX),
		.CurrentY(CurrentY),
		.mapData(hallwayTop),
		.wall(playerColor)
	);
	
	HallwayRight HallwayRight(
		.clk_vga(clk_vga),
		.CurrentX(CurrentX),
		.CurrentY(CurrentY),
		.mapData(hallwayRight),
		.wall(playerColor)
	);
	
	BlackKeyRoom BlackKeyRoom(
		.clk_vga(clk_vga),
		.CurrentX(CurrentX),
		.CurrentY(CurrentY),
		.mapData(blackKeyRoom),
		.wall(playerColor)
	);
	
	HallwayLeft HallwayLeft(
		.clk_vga(clk_vga),
		.CurrentX(CurrentX),
		.CurrentY(CurrentY),
		.mapData(hallwayLeft),
		.wall(playerColor)
	);
	
	
	
	//Draws the map based on the current mapX and mapY
	//The idea is to have only one output from the map generator module
	//And do all the heavy lifting in the top module
	//The map generator acts as a datapath for the static objects in the game
	always @(posedge clk_vga) begin
		if(HBlank || VBlank) begin
			mColor <= 0;
		end
		else begin
			
			//VGA test pattern for debugging purposes
			/*
			if(CurrentY < 160) begin
				mColor[7:5] <= 3'b111;
			end
			else if(CurrentY < 320) begin
				mColor[4:2] <= 3'b111;
			end
			else begin
				mColor[1:0] <= 2'b11;
			end
			*/
				
			//Starting castle
			if(mapX == 3 && mapY == 5) begin
				mColor[7:0] <= startCastle[7:0];
			end 
			//Central hallway
			else if(mapX == 3 && mapY == 6) begin
				mColor[7:0] <= hallwayTop[7:0];
			end 
			//Right hallway
			else if(mapX == 4 && mapY == 6) begin
				mColor[7:0] <= hallwayRight[7:0];
			end
			//Black key room
			else if(mapX == 4 && mapY == 7) begin
				mColor[7:0] <= blackKeyRoom[7:0];
			end
			//Left hallway
			else if(mapX == 2 && mapY == 6) begin
				mColor[7:0] <= hallwayLeft;
			end
			else begin
				mColor[7:0] <= 8'b00000000;
			end
			
		end
	end
	
	assign mapData[7:0] = mColor[7:0];
	
endmodule
